`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/07/2017 10:23:29 AM
// Design Name: 
// Module Name: Datapath
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module Datapath();

reg clk;
//Clock initialization
initial
begin
    clk = 0;
    forever #25 clk = ~clk;
end

wire exempt_zero, exempt_neg;
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// IF Section Wires
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire [31:0] pc_in;
wire [31:0] pc_out; 
wire [31:0] pc_plus1;
wire [31:0] im_out;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//ID Section Wires
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire [31:0] rs_out, rt_out;
wire [31:0] id_out;
wire [31:0] sign_out;
wire [31:0] id_alu;
wire [31:0] ext_alu;
wire RegWrt, MemToReg, PCToReg, BranchNeg, BranchZero, Jump, JumpMem, MemRead, MemWrt;
wire [3:0] ALUOp;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//EX Section Wires
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire ex_RegWrt, ex_MemToReg, ex_PCToReg, ex_BranchNeg, ex_BranchZero, ex_Jump, ex_JumpMem, ex_MemRead, ex_MemWrt, ex_N, ex_Z;
wire [31:0] ex_rs, ex_rt, ex_data_out, ex_ext_alu, ex_alu;
wire [5:0] ex_rd;
wire [3:0] ex_ALUOP;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//WB Section Wires
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

wire wb_RegWrt, wb_MemToReg, wb_PCToReg, wb_BranchNeg, wb_BranchZero, wb_Jump, wb_JumpMem, wb_N, wb_Z;
wire controlA, controlB, Branch_result;
wire [31:0] wb_alu, wb_data_out, wb_mux, wb_ext_alu;
wire [5:0] wb_rd;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
// Datapath 
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////


///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//IF Section
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//Calling Mux before PC
ThreeToOne PCMux(controlA, controlB, pc_plus1, wb_alu, wb_data_out );

//Program Counter 
PC prog_counter(clk, pc_plus1, pc_out); 

//Increment PC by 1
ArithmeticLogicUnit IncrementPC(pc_out, pc_out, 4'b0001, pc_plus1, exempt_zero, exempt_neg);

//Instruction Memory
InstructionMemory InstrMem(pc_out, clk, im_out);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//ID Section
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//IF_ID buffer
IF_ID_Buf IFIDBuf(clk, im_out, id_out, pc_out, id_alu);

//COntrol
Control idControl( clk, id_out[31:28], RegWrt, MemToReg, PCToReg, BranchNeg, BranchZero, Jump, JumpMem, ALUOp, MemRead, MemWrt);

//Register Memory
wire [5:0] test_RM_rs, test_RM_rt, test_RM_rd;
RegisterMemory RegMemory(id_out[21:16], id_out[15:10], id_out[27:22], wb_mux, wb_RegWrt, rs_out, rt_out, clk, test_RM_rs, test_RM_rt, test_RM_rd);

//Sign Extend
SignExtend extend(clk, id_out[21:0], sign_out);

//ID ALU
ArithmeticLogicUnit idALU(sign_out, id_alu, 4'b0000, ext_alu, exempt_zero, exempt_neg);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//EX Sections
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//ID_EX Buffer
ID_EX_Buf IDEXBuf(clk, RegWrt, MemToReg, PCToReg, BranchNeg, ALUOp, MemRead, MemWrt,BranchZero, Jump, JumpMem, rs_out, rt_out, id_out[27:22], sign_out, 
                     ex_RegWrt, ex_MemToReg, ex_PCToReg, ex_BranchNeg, ex_ALUOP, ex_MemRead, ex_MemWrt,ex_BranchZero, ex_Jump, ex_JumpMem, ex_rs, ex_rt, ex_rd, ex_ext_alu );

//Data Memory
DataMemory D_memory(clk, ex_MemWrt, ex_MemRead, ex_rs, ex_rt, ex_data_out);

//EX ALU
wire [31:0] testA, testB, testOpcode, testResult, testInternalA;
ArithmeticLogicUnit exALU(ex_rs, ex_rt,ex_ALUOP, ex_alu, ex_Z, ex_N, testA, testB, testInternalA, testOpcode, testResult);

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
//WB Section
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

//EX_WB Buffer
 EX_WB_Buf exwBuf(clk, ex_N, ex_Z, ex_RegWrt,ex_MemToReg, ex_PCToReg, ex_BranchNeg, ex_BranchZero, ex_Jump, ex_JumpMem, ex_alu, ex_data_out, ex_rd, ex_ext_alu,
                     wb_N, wb_Z, wb_RegWrt,wb_MemToReg, wb_PCToReg, wb_BranchNeg, wb_BranchZero, wb_Jump, wb_JumpMem, wb_alu, wb_data_out, wb_rd, wb_ext_alu);

//WB Mux
ThreeToOne wbMux(wb_PCToReg, wb_MemToReg, wb_alu, wb_data_out, wb_ext_alu, wb_mux);

//PCSource to get control for IF Mux
PCSource branch(ex_N, ex_Z, ex_BranchNeg, ex_BranchZero, ex_Jump, ex_JumpMem, controlA, controlB);


endmodule
